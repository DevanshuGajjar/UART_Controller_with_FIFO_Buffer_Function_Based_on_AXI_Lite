`timescale 1ns/1ps


module BAUDGEN
(
	input			clk,
	input			a_resetn,
	input		[3:0]	baudrate,

	output	reg		baudtick
);



endmodule

